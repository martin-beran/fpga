-- Demo of library package lib_io.pkg_vga

library ieee;
use ieee.std_logic_1164.all;

entity demo_vga is
	port (
	);
end entity;

architecture main of demo_vga is
begin
end architecture;