-- MB50: CDI (Control and Debugging Interface)

entity cdi is
	port (
	);
end entity;

architecture main of cdi is
begin
end architecture;