-- MB50 main entity, it composes all components of computer MB50

entity mb50 is
begin
end entity;

architecture main of mb50 is
begin
end architecture;