-- Clock adapters

library ieee;
use ieee.std_logic_1164.all;

package pkg_clock is
	-- Divider of an input clock frequency.
	-- Generates pulses of a length equal to the period of the master clock at
	-- some rising edges of the input clock.
	component clock_divider is
		generic (
			-- number of input clock periods between output pulses
			factor: positive range 2 to positive'high
		);
		port (
			-- the master system clock
			Clk: in std_logic;
			-- Reset and start from the beginning
			Rst: in std_logic := '0';
			-- the input synchronization from a previous level clock_divider
			ISync: in std_logic := '1';
			-- the output clock (registered)
			O: out std_logic;
			-- the output synchronization signal for a next level clock_subdivider (unregistered)
			OSync: out std_logic
		);
	end component;
	
	-- Toggle the output with each input pulse
	-- It converts pulses generated by clock_divider to a signal with duty cycle 50 % with
	-- half frequency
	component half_f_duty_50 is
		port (
			-- the master system clock
			Clk: in std_logic;
			-- Reset and start from the beginning
			Rst: in std_logic;
			-- the input clock (expected
			I: in std_logic;
			-- the output signal
			O: out std_logic
		);
	end component;
end package;

-- clock divider --------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library lib_util;
use lib_util.pkg_clock.all;

entity clock_divider is
	generic (
		factor: positive
	);
	port (
		Clk, Rst, ISync: in std_logic;
		O, OSync: out std_logic
	);
end entity;

architecture main of clock_divider is
	signal f: natural range 0 to factor - 1 := factor - 1;
begin
	OSync <= ISync when f = factor - 1 else '0';
	process (Clk, Rst) is
	begin
		if Rst then
			f <= factor - 1;
			O <= '0';
		elsif rising_edge(Clk) then
			O <= '0';
			if ISync = '1' then
				if f = factor - 1 then
					f <= 0;
					O <= '1';
				else
					f <= f + 1;
				end if;
			end if;
		end if;
	end process;
end architecture;

-- half_f_duty_50 -------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library lib_util;
use lib_util.pkg_clock.all;

entity half_f_duty_50 is
	port (
		Clk, Rst, I: in std_logic;
		O: out std_logic
	);
end entity;

architecture main of half_f_duty_50 is
begin
	process (Clk, Rst, I) is
	begin
		if rising_edge(Clk) then
			if Rst = '1' then
				O <= '0';
			elsif I = '1' then
				O <= not O;
			end if;
		end if;
	end process;
end architecture;