-- VGA controller

library ieee;
use ieee.std_logic_1164;

package pkg_vga is
	component vga is
		port (
		);
	end component;
end package;

library ieee;
use ieee.std_logic_1164;

entity vga is
	port (
	);
end entity;

architecture main of vga is
begin
end architecture;