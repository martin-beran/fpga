-- Time keeping

library ieee;
use ieee.std_logic_1164.all;

entity counter is
	generic (
		-- TODO
	);
	port (
		-- TODO
	);
end entity;

architecture main of counter is
begin
	-- TODO
end architecture;