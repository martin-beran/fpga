-- Demo of library package lib_io.pkg_uart

library ieee;
use ieee.std_logic_1164.all;

entity demo_uart is
	port (
	);
end entity;

architecture main of demo_uart is
begin
end architecture;