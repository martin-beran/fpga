-- Parameters of the system master clock crystal

package pkg_crystal is
	-- Frequency of the system master clock crystal
	constant crystal_hz: positive := 50_000_000;
end package;